LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY data_in IS
	GENERIC(DATA_WIDTH: INTEGER;
		ROW_SIZE: INTEGER;
		COL_SIZE: INTEGER);
	PORT(	Clk: IN STD_LOGIC;
		We_in: IN STD_LOGIC;
		Re_in: IN STD_LOGIC;
		Addr: IN INTEGER RANGE 0 TO COL_SIZE * ROW_SIZE - 1;
		Data_in: IN INTEGER RANGE 0 TO 2**DATA_WIDTH - 1;
		Data_out: OUT INTEGER RANGE 0 TO 2**DATA_WIDTH - 1);
END data_in;

ARCHITECTURE data_in_arch OF data_in IS
	TYPE DATA_ARRAY IS ARRAY(0 TO COL_SIZE * ROW_SIZE - 1) OF INTEGER;
	SIGNAL Matrix_in : DATA_ARRAY := (62, 124, 129, 129, 190, 221, 88, 138, 217, 205, 186, 14, 217, 215, 253, 37, 220, 50, 97, 54, 235, 171, 69, 246, 210, 17, 178, 240, 135, 174, 97, 169,
3, 159, 77, 131, 39, 45, 19, 199, 218, 204, 210, 28, 175, 195, 220, 22, 126, 61, 237, 101, 74, 203, 84, 148, 117, 213, 29, 125, 91, 155, 26, 150,
227, 49, 175, 201, 90, 135, 127, 148, 75, 190, 108, 252, 137, 40, 177, 222, 15, 49, 189, 37, 247, 73, 53, 197, 43, 87, 216, 104, 149, 181, 159, 211,
59, 210, 35, 72, 73, 8, 230, 199, 68, 60, 36, 113, 245, 48, 234, 236, 30, 142, 163, 236, 7, 18, 21, 249, 248, 83, 129, 57, 1, 18, 225, 20,
42, 152, 247, 103, 13, 240, 130, 195, 252, 120, 52, 150, 174, 8, 211, 122, 12, 4, 189, 48, 4, 201, 13, 86, 39, 124, 6, 21, 133, 224, 164, 29,
142, 213, 134, 208, 208, 223, 235, 51, 170, 231, 238, 73, 88, 9, 161, 126, 56, 56, 239, 71, 72, 181, 155, 224, 165, 224, 68, 200, 123, 191, 123, 20,
28, 203, 135, 100, 113, 49, 10, 16, 164, 69, 232, 188, 224, 6, 137, 163, 106, 58, 29, 115, 206, 213, 212, 72, 47, 62, 10, 35, 59, 16, 47, 124,
61, 10, 101, 48, 79, 243, 200, 117, 11, 29, 140, 78, 74, 184, 88, 122, 99, 189, 131, 198, 87, 103, 72, 63, 221, 157, 207, 213, 179, 170, 63, 181,
209, 40, 100, 56, 67, 61, 161, 155, 126, 46, 38, 34, 12, 72, 251, 244, 44, 109, 153, 190, 70, 204, 230, 203, 188, 202, 77, 224, 110, 127, 153, 102,
114, 88, 133, 169, 153, 44, 202, 32, 7, 129, 253, 84, 143, 243, 234, 252, 246, 231, 224, 19, 248, 3, 219, 2, 74, 233, 240, 188, 194, 210, 2, 32,
163, 58, 2, 215, 138, 67, 67, 235, 210, 26, 78, 79, 135, 26, 245, 31, 123, 203, 194, 175, 134, 134, 244, 52, 200, 181, 109, 36, 226, 105, 75, 113,
117, 249, 184, 246, 139, 191, 32, 169, 44, 175, 11, 144, 30, 43, 5, 180, 116, 244, 211, 201, 71, 225, 70, 69, 229, 139, 253, 82, 223, 118, 251, 179,
118, 30, 43, 15, 91, 55, 218, 231, 98, 123, 152, 148, 250, 177, 173, 35, 201, 121, 164, 213, 60, 96, 74, 95, 51, 161, 21, 144, 149, 113, 168, 141,
189, 67, 114, 133, 109, 149, 81, 217, 206, 76, 46, 124, 19, 45, 161, 178, 229, 221, 149, 232, 64, 40, 166, 23, 252, 106, 170, 151, 133, 171, 89, 127,
87, 46, 12, 92, 170, 218, 103, 203, 4, 132, 146, 52, 220, 48, 214, 199, 180, 163, 54, 152, 177, 206, 181, 164, 40, 45, 230, 199, 84, 231, 238, 76,
150, 135, 93, 129, 22, 203, 176, 5, 19, 31, 91, 58, 196, 147, 107, 226, 45, 58, 248, 0, 118, 151, 41, 150, 75, 145, 32, 77, 126, 225, 190, 86,
88, 37, 147, 202, 207, 193, 111, 165, 246, 4, 94, 36, 25, 30, 200, 48, 53, 99, 147, 37, 91, 74, 119, 115, 235, 164, 96, 160, 211, 211, 155, 73,
230, 87, 212, 168, 132, 196, 214, 137, 250, 117, 25, 193, 68, 248, 64, 98, 58, 208, 100, 239, 154, 222, 18, 169, 67, 42, 157, 99, 88, 92, 69, 150,
213, 235, 48, 239, 20, 55, 162, 93, 230, 165, 169, 78, 215, 53, 178, 50, 152, 160, 169, 80, 79, 124, 242, 82, 142, 190, 42, 204, 140, 11, 57, 184,
22, 101, 251, 95, 62, 29, 69, 242, 28, 30, 240, 115, 246, 101, 76, 225, 139, 44, 49, 127, 112, 148, 32, 125, 221, 137, 227, 191, 230, 170, 163, 35,
103, 229, 22, 22, 198, 223, 48, 123, 5, 54, 199, 28, 214, 141, 52, 102, 139, 63, 209, 4, 233, 210, 211, 86, 17, 131, 188, 25, 72, 107, 70, 37,
226, 101, 101, 90, 26, 128, 250, 163, 251, 117, 100, 7, 228, 244, 19, 156, 86, 117, 105, 177, 166, 21, 65, 142, 209, 23, 2, 251, 121, 159, 102, 54,
108, 250, 10, 85, 110, 20, 39, 2, 52, 156, 240, 218, 176, 18, 236, 44, 153, 222, 174, 37, 114, 22, 178, 70, 72, 213, 167, 253, 166, 24, 10, 105,
85, 223, 84, 36, 216, 8, 26, 17, 34, 19, 230, 125, 248, 24, 46, 116, 235, 171, 130, 92, 91, 49, 167, 106, 176, 191, 179, 174, 203, 150, 173, 178,
228, 179, 17, 31, 85, 95, 29, 138, 103, 102, 146, 55, 144, 38, 231, 73, 17, 177, 22, 93, 245, 67, 108, 37, 33, 247, 253, 132, 68, 70, 165, 157,
102, 223, 209, 49, 176, 22, 232, 188, 148, 191, 106, 91, 30, 222, 8, 91, 67, 189, 75, 164, 254, 38, 58, 144, 40, 38, 194, 241, 176, 235, 65, 154,
181, 165, 140, 117, 45, 125, 101, 73, 13, 197, 17, 84, 6, 62, 113, 148, 125, 120, 107, 221, 46, 145, 192, 26, 214, 106, 3, 148, 109, 44, 206, 169,
125, 5, 146, 60, 187, 150, 196, 146, 172, 222, 101, 108, 162, 252, 46, 3, 235, 167, 126, 122, 18, 225, 199, 25, 29, 119, 136, 103, 114, 178, 214, 189,
222, 12, 153, 24, 108, 162, 56, 182, 177, 195, 182, 239, 146, 204, 207, 143, 109, 121, 52, 38, 89, 109, 7, 101, 94, 154, 191, 202, 42, 138, 186, 173,
246, 247, 33, 180, 102, 43, 77, 128, 242, 143, 237, 202, 101, 17, 92, 144, 183, 124, 126, 252, 22, 208, 41, 201, 183, 17, 66, 196, 192, 139, 21, 36,
187, 245, 217, 40, 58, 231, 254, 180, 206, 102, 112, 88, 141, 40, 194, 79, 146, 219, 162, 193, 97, 184, 193, 214, 22, 157, 240, 205, 102, 47, 241, 131,
42, 71, 214, 222, 14, 93, 77, 188, 156, 4, 73, 217, 30, 166, 248, 56, 135, 175, 133, 29, 55, 236, 143, 10, 196, 230, 99, 140, 194, 233, 167, 219
);
	BEGIN
		PROCESS(Clk)
		BEGIN
			IF (Clk'Event AND Clk = '1') THEN
				IF (We_in = '1') THEN Matrix_in(Addr) <= Data_in;
				ELSE 
					IF (Re_in = '1') THEN Data_out <= Matrix_in(Addr);
					END IF;
				END IF;
			END IF;
		END PROCESS;
END data_in_arch;
