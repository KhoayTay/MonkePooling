LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE my_package IS

COMPONENT counter IS
	GENERIC(stop_value: INTEGER);
	PORT(	Clk, Inc, Clr: IN STD_LOGIC;
		Z: OUT STD_LOGIC;
		Count: OUT INTEGER RANGE 0 TO stop_value);
END COMPONENT;

COMPONENT data_in IS
	GENERIC(DATA_WIDTH: INTEGER;
		ROW_SIZE: INTEGER;
		COL_SIZE: INTEGER);
	PORT(	Clk: IN STD_LOGIC;
		We_in: IN STD_LOGIC;
		Re_in: IN STD_LOGIC;
		Addr: IN INTEGER RANGE 0 TO ROW_SIZE * COL_SIZE - 1;
		Data_in: IN INTEGER RANGE 0 TO 2**DATA_WIDTH - 1;
		Data_out: OUT INTEGER RANGE 0 TO 2**DATA_WIDTH - 1);		
END COMPONENT;

COMPONENT data_out IS
	GENERIC(DATA_WIDTH: INTEGER;
		ROW_SIZE: INTEGER;
		COL_SIZE: INTEGER);
	PORT(	Clk: IN STD_LOGIC;
		We_out: IN STD_LOGIC;
		Re_out: IN STD_LOGIC;
		Clean: IN STD_LOGIC;
		Addr: IN INTEGER RANGE 0 TO COL_SIZE * ROW_SIZE - 1;
		Data_in: IN INTEGER RANGE 0 TO 2**DATA_WIDTH - 1;
		Data_out: OUT INTEGER RANGE 0 TO 2**DATA_WIDTH - 1;
		Done: OUT STD_LOGIC);		
END COMPONENT;

COMPONENT datapath IS
	GENERIC(DATA_WIDTH: INTEGER;
		ROW_SIZE_IN: INTEGER;
		COL_SIZE_IN: INTEGER;
		ROW_SIZE_OUT: INTEGER;
		COL_SIZE_OUT: INTEGER;
		ROW_STEP: INTEGER;
		COL_STEP: INTEGER);
	PORT(	Clk: IN STD_LOGIC;
		R_clr, Rs_clr, C_clr, Cs_clr: IN STD_LOGIC;
		R_inc, Rs_inc, C_inc, Cs_inc: IN STD_LOGIC;
		Data_in, Data_out: IN INTEGER RANGE 0 TO 2**DATA_WIDTH - 1;
		R_z, Rs_z, C_z, Cs_z: OUT STD_LOGIC;
		Data_in_addr: OUT INTEGER RANGE 0 TO ROW_SIZE_IN * COL_SIZE_IN - 1;
		Data_out_addr: OUT INTEGER RANGE 0 TO ROW_SIZE_OUT * COL_SIZE_OUT - 1;
		New_data_out: OUT INTEGER RANGE 0 TO 2**DATA_WIDTH - 1);
END COMPONENT;

COMPONENT controller IS
	GENERIC(DATA_WIDTH: INTEGER);
	PORT(	Start: IN STD_LOGIC;
		Clk: IN STD_LOGIC;
		Reset: IN STD_LOGIC;
		Done_Clean: IN STD_LOGIC;
		R_z, Rs_z, C_z, Cs_z: IN STD_LOGIC;
		R_clr, Rs_Clr, C_clr, Cs_clr: OUT STD_LOGIC;
		R_inc, Rs_inc, C_inc, Cs_inc: OUT STD_LOGIC;
		Re_in, Re_out, We_in, We_out: OUT STD_LOGIC;
		Clean: OUT STD_LOGIC;
		Done: OUT STD_LOGIC);
END COMPONENT;

COMPONENT pooling IS
	GENERIC(DATA_WIDTH: INTEGER;
		ROW_SIZE_IN: INTEGER;
		COL_SIZE_IN: INTEGER;
		ROW_SIZE_OUT: INTEGER;
		COL_SIZE_OUT: INTEGER;
		ROW_STEP: INTEGER;
		COL_STEP: INTEGER);
	PORT(	Clk: IN STD_LOGIC;
		Start: IN STD_LOGIC;
		Reset: IN STD_LOGIC;		
		Done: OUT STD_LOGIC);	
END COMPONENT;	

END PACKAGE my_package;
